module psi

pub struct LineComment {
	PsiElementImpl
}

pub struct BlockComment {
	PsiElementImpl
}
